library verilog;
use verilog.vl_types.all;
entity maq_estado_vlg_vec_tst is
end maq_estado_vlg_vec_tst;
