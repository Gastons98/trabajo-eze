library verilog;
use verilog.vl_types.all;
entity maq_estado_vlg_check_tst is
    port(
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        d4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end maq_estado_vlg_check_tst;
