library verilog;
use verilog.vl_types.all;
entity ej_combinacional_vlg_check_tst is
    port(
        led             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ej_combinacional_vlg_check_tst;
