library verilog;
use verilog.vl_types.all;
entity sumador_completo_vlg_check_tst is
    port(
        coutsuma        : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end sumador_completo_vlg_check_tst;
