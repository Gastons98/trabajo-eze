library verilog;
use verilog.vl_types.all;
entity ej_combinacional_vlg_vec_tst is
end ej_combinacional_vlg_vec_tst;
