library verilog;
use verilog.vl_types.all;
entity sumador_completo_ffD_vlg_check_tst is
    port(
        out_cout        : in     vl_logic;
        out_suma        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sumador_completo_ffD_vlg_check_tst;
